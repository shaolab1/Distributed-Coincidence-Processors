parameter int DELAY_PAIR = 104;
parameter int CHAN_DELAY_MAT[PAIR_NUM][2] = '{'{4,1},'{4,2},'{4,0},'{4,1},'{4,5},'{4,5},'{4,3},'{4,0},'{4,1},'{4,2},'{4,4},'{4,0},'{4,0},
                                              '{2,2},'{2,0},'{2,1},'{2,5},'{2,5},'{2,3},'{2,0},'{2,1},'{2,2},'{2,4},'{2,0},'{2,0},'{2,1},
                                              '{1,0},'{1,1},'{1,5},'{1,5},'{1,3},'{1,0},'{1,1},'{1,2},'{1,4},'{1,0},'{1,0},'{1,1},
                                              '{2,1},'{2,5},'{2,5},'{2,3},'{2,0},'{2,1},'{2,2},'{2,4},'{2,0},'{2,0},'{2,1},
                                              '{0,5},'{0,5},'{0,3},'{0,0},'{0,1},'{0,2},'{0,4},'{0,0},'{0,0},'{0,1},
                                              '{1,5},'{1,3},'{1,0},'{1,1},'{1,2},'{1,4},'{1,0},'{1,0},'{1,1},
                                              '{5,3},'{5,0},'{5,1},'{5,2},'{5,4},'{5,0},'{5,0},'{5,1},
                                              '{5,0},'{5,1},'{5,2},'{5,4},'{5,0},'{5,0},'{5,1},
                                              '{3,1},'{3,2},'{3,4},'{3,0},'{3,0},'{3,1},
                                              '{0,2},'{0,4},'{0,0},'{0,0},'{0,1},
                                              '{1,4},'{1,0},'{1,0},'{1,1},
                                              '{2,0},'{2,0},'{2,1},
                                              '{4,0},'{4,1},
                                              '{0,1}};